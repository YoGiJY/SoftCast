
`resetall
`timescale 1ns/1ps
module ROM5_omega (ROM_data, ROM_addr,clk);
  
  parameter WORDLENGTH=18,ADDRLENGTH=10;
  
  output [WORDLENGTH-1:0] ROM_data;
  input 	[ADDRLENGTH-1:0] ROM_addr;
  input  clk;
  reg    [WORDLENGTH-1:0] ROM_data;
  
  always @ (posedge clk)
  begin
    case(ROM_addr)
        10'b0000000000:ROM_data<=18'b011111111000000000;
        10'b0000000001:ROM_data<=18'b011111111000000000;
        10'b0000000010:ROM_data<=18'b011111111000000000;
        10'b0000000011:ROM_data<=18'b011111111000000000;
        10'b0000000100:ROM_data<=18'b011111111000000000;
        10'b0000000101:ROM_data<=18'b011101011110011111;
        10'b0000000110:ROM_data<=18'b010110100101001100;
        10'b0000000111:ROM_data<=18'b001100001100010101;
        10'b0000001000:ROM_data<=18'b011111111000000000;
        10'b0000001001:ROM_data<=18'b010110100101001100;
        10'b0000001010:ROM_data<=18'b000000000100000001;
        10'b0000001011:ROM_data<=18'b101001100101001100;
        10'b0000001100:ROM_data<=18'b011111111000000000;
        10'b0000001101:ROM_data<=18'b001100001100010101;
        10'b0000001110:ROM_data<=18'b101001100101001100;
        10'b0000001111:ROM_data<=18'b100010101001100001;
        10'b0000010000:ROM_data<=18'b011111111000000000;
        10'b0000010001:ROM_data<=18'b011111101111101000;
        10'b0000010010:ROM_data<=18'b011111010111001111;
        10'b0000010011:ROM_data<=18'b011110100110110110;
        10'b0000010100:ROM_data<=18'b011111111000000000;
        10'b0000010101:ROM_data<=18'b011100000110001000;
        10'b0000010110:ROM_data<=18'b010001101100101100;
        10'b0000010111:ROM_data<=18'b000011000100000011;
        10'b0000011000:ROM_data<=18'b011111111000000000;
        10'b0000011001:ROM_data<=18'b010100001100111011;
        10'b0000011010:ROM_data<=18'b111001111100000110;
        10'b0000011011:ROM_data<=18'b100100000110001000;
        10'b0000011100:ROM_data<=18'b011111111000000000;
        10'b0000011101:ROM_data<=18'b001001010100001100;
        10'b0000011110:ROM_data<=18'b100101100101110011;
        10'b0000011111:ROM_data<=18'b100111011010100001;
        10'b0000100000:ROM_data<=18'b011111111000000000;
        10'b0000100001:ROM_data<=18'b011111010111001111;
        10'b0000100010:ROM_data<=18'b011101011110011111;
        10'b0000100011:ROM_data<=18'b011010100101110011;
        10'b0000100100:ROM_data<=18'b011111111000000000;
        10'b0000100101:ROM_data<=18'b011010100101110011;
        10'b0000100110:ROM_data<=18'b001100001100010101;
        10'b0000100111:ROM_data<=18'b111001111100000110;
        10'b0000101000:ROM_data<=18'b011111111000000000;
        10'b0000101001:ROM_data<=18'b010001101100101100;
        10'b0000101010:ROM_data<=18'b110011111100010101;
        10'b0000101011:ROM_data<=18'b100000110111001111;
        10'b0000101100:ROM_data<=18'b011111111000000000;
        10'b0000101101:ROM_data<=18'b000110001100000110;
        10'b0000101110:ROM_data<=18'b100010101110011111;
        10'b0000101111:ROM_data<=18'b101110011011010100;
        10'b0000110000:ROM_data<=18'b011111111000000000;
        10'b0000110001:ROM_data<=18'b011110100110110110;
        10'b0000110010:ROM_data<=18'b011010100101110011;
        10'b0000110011:ROM_data<=18'b010100001100111011;
        10'b0000110100:ROM_data<=18'b011111111000000000;
        10'b0000110101:ROM_data<=18'b011000101101011111;
        10'b0000110110:ROM_data<=18'b000110001100000110;
        10'b0000110111:ROM_data<=18'b110001000100100000;
        10'b0000111000:ROM_data<=18'b011111111000000000;
        10'b0000111001:ROM_data<=18'b001111000100100000;
        10'b0000111010:ROM_data<=18'b101110011100101100;
        10'b0000111011:ROM_data<=18'b100000011000011000;
        10'b0000111100:ROM_data<=18'b011111111000000000;
        10'b0000111101:ROM_data<=18'b000011000100000011;
        10'b0000111110:ROM_data<=18'b100000110111001111;
        10'b0000111111:ROM_data<=18'b110110110011110100;
        10'b0001000000:ROM_data<=18'b011111111000000000;
        10'b0001000001:ROM_data<=18'b011111110111111010;
        10'b0001000010:ROM_data<=18'b011111110111110100;
        10'b0001000011:ROM_data<=18'b011111110111101110;
        10'b0001000100:ROM_data<=18'b011111111000000000;
        10'b0001000101:ROM_data<=18'b011101001110011001;
        10'b0001000110:ROM_data<=18'b010101011101000100;
        10'b0001000111:ROM_data<=18'b001001111100001110;
        10'b0001001000:ROM_data<=18'b011111111000000000;
        10'b0001001001:ROM_data<=18'b010101111101001000;
        10'b0001001010:ROM_data<=18'b111110100100000010;
        10'b0001001011:ROM_data<=18'b100111111101011010;
        10'b0001001100:ROM_data<=18'b011111111000000000;
        10'b0001001101:ROM_data<=18'b001011011100010011;
        10'b0001001110:ROM_data<=18'b101000100101010101;
        10'b0001001111:ROM_data<=18'b100011101001110010;
        10'b0001010000:ROM_data<=18'b011111111000000000;
        10'b0001010001:ROM_data<=18'b011111101111100001;
        10'b0001010010:ROM_data<=18'b011110111111000011;
        10'b0001010011:ROM_data<=18'b011101101110100101;
        10'b0001010100:ROM_data<=18'b011111111000000000;
        10'b0001010101:ROM_data<=18'b011011101110000011;
        10'b0001010110:ROM_data<=18'b010000011100100110;
        10'b0001010111:ROM_data<=18'b000000110100000010;
        10'b0001011000:ROM_data<=18'b011111111000000000;
        10'b0001011001:ROM_data<=18'b010011100100110111;
        10'b0001011010:ROM_data<=18'b111000011100001001;
        10'b0001011011:ROM_data<=18'b100010111110011001;
        10'b0001011100:ROM_data<=18'b011111111000000000;
        10'b0001011101:ROM_data<=18'b001000100100001011;
        10'b0001011110:ROM_data<=18'b100100110101111101;
        10'b0001011111:ROM_data<=18'b101001000010101111;
        10'b0001100000:ROM_data<=18'b011111111000000000;
        10'b0001100001:ROM_data<=18'b011111000111001001;
        10'b0001100010:ROM_data<=18'b011100110110010011;
        10'b0001100011:ROM_data<=18'b011001001101100100;
        10'b0001100100:ROM_data<=18'b011111111000000000;
        10'b0001100101:ROM_data<=18'b011010000101101110;
        10'b0001100110:ROM_data<=18'b001010101100010000;
        10'b0001100111:ROM_data<=18'b110111100100001011;
        10'b0001101000:ROM_data<=18'b011111111000000000;
        10'b0001101001:ROM_data<=18'b010001000100101001;
        10'b0001101010:ROM_data<=18'b110010011100011010;
        10'b0001101011:ROM_data<=18'b100000011111100001;
        10'b0001101100:ROM_data<=18'b011111111000000000;
        10'b0001101101:ROM_data<=18'b000101011100000101;
        10'b0001101110:ROM_data<=18'b100010000110101011;
        10'b0001101111:ROM_data<=18'b110000011011011101;
        10'b0001110000:ROM_data<=18'b011111111000000000;
        10'b0001110001:ROM_data<=18'b011110010110110001;
        10'b0001110010:ROM_data<=18'b011001100101101001;
        10'b0001110011:ROM_data<=18'b010010010100110000;
        10'b0001110100:ROM_data<=18'b011111111000000000;
        10'b0001110101:ROM_data<=18'b011000001101011010;
        10'b0001110110:ROM_data<=18'b000100101100000100;
        10'b0001110111:ROM_data<=18'b101111000100101001;
        10'b0001111000:ROM_data<=18'b011111111000000000;
        10'b0001111001:ROM_data<=18'b001110010100011101;
        10'b0001111010:ROM_data<=18'b101101001100110100;
        10'b0001111011:ROM_data<=18'b100000101000101011;
        10'b0001111100:ROM_data<=18'b011111111000000000;
        10'b0001111101:ROM_data<=18'b000010010100000010;
        10'b0001111110:ROM_data<=18'b100000100111011011;
        10'b0001111111:ROM_data<=18'b111001001011111000;
        10'b0010000000:ROM_data<=18'b011111111000000000;
        10'b0010000001:ROM_data<=18'b011111110111110100;
        10'b0010000010:ROM_data<=18'b011111101111101000;
        10'b0010000011:ROM_data<=18'b011111100111011011;
        10'b0010000100:ROM_data<=18'b011111111000000000;
        10'b0010000101:ROM_data<=18'b011100110110010011;
        10'b0010000110:ROM_data<=18'b010100001100111011;
        10'b0010000111:ROM_data<=18'b000111101100001001;
        10'b0010001000:ROM_data<=18'b011111111000000000;
        10'b0010001001:ROM_data<=18'b010101011101000100;
        10'b0010001010:ROM_data<=18'b111101000100000011;
        10'b0010001011:ROM_data<=18'b100110100101101001;
        10'b0010001100:ROM_data<=18'b011111111000000000;
        10'b0010001101:ROM_data<=18'b001010101100010000;
        10'b0010001110:ROM_data<=18'b100111011101011111;
        10'b0010001111:ROM_data<=18'b100100110010000011;
        10'b0010010000:ROM_data<=18'b011111111000000000;
        10'b0010010001:ROM_data<=18'b011111100111011011;
        10'b0010010010:ROM_data<=18'b011110100110110110;
        10'b0010010011:ROM_data<=18'b011100110110010011;
        10'b0010010100:ROM_data<=18'b011111111000000000;
        10'b0010010101:ROM_data<=18'b011011010101111101;
        10'b0010010110:ROM_data<=18'b001111000100100000;
        10'b0010010111:ROM_data<=18'b111110100100000010;
        10'b0010011000:ROM_data<=18'b011111111000000000;
        10'b0010011001:ROM_data<=18'b010010111100110100;
        10'b0010011010:ROM_data<=18'b110110110100001100;
        10'b0010011011:ROM_data<=18'b100010000110101011;
        10'b0010011100:ROM_data<=18'b011111111000000000;
        10'b0010011101:ROM_data<=18'b000111101100001001;
        10'b0010011110:ROM_data<=18'b100100000110001000;
        10'b0010011111:ROM_data<=18'b101010101010111100;
        10'b0010100000:ROM_data<=18'b011111111000000000;
        10'b0010100001:ROM_data<=18'b011110111111000011;
        10'b0010100010:ROM_data<=18'b011100000110001000;
        10'b0010100011:ROM_data<=18'b010111100101010101;
        10'b0010100100:ROM_data<=18'b011111111000000000;
        10'b0010100101:ROM_data<=18'b011001100101101001;
        10'b0010100110:ROM_data<=18'b001001010100001100;
        10'b0010100111:ROM_data<=18'b110101011100010000;
        10'b0010101000:ROM_data<=18'b011111111000000000;
        10'b0010101001:ROM_data<=18'b010000011100100110;
        10'b0010101010:ROM_data<=18'b110001000100100000;
        10'b0010101011:ROM_data<=18'b100000010111110100;
        10'b0010101100:ROM_data<=18'b011111111000000000;
        10'b0010101101:ROM_data<=18'b000100101100000100;
        10'b0010101110:ROM_data<=18'b100001100110110110;
        10'b0010101111:ROM_data<=18'b110010011011100110;
        10'b0010110000:ROM_data<=18'b011111111000000000;
        10'b0010110001:ROM_data<=18'b011110000110101011;
        10'b0010110010:ROM_data<=18'b011000101101011111;
        10'b0010110011:ROM_data<=18'b010000011100100110;
        10'b0010110100:ROM_data<=18'b011111111000000000;
        10'b0010110101:ROM_data<=18'b010111100101010101;
        10'b0010110110:ROM_data<=18'b000011000100000011;
        10'b0010110111:ROM_data<=18'b101101001100110100;
        10'b0010111000:ROM_data<=18'b011111111000000000;
        10'b0010111001:ROM_data<=18'b001101101100011010;
        10'b0010111010:ROM_data<=18'b101011111100111011;
        10'b0010111011:ROM_data<=18'b100001001000111101;
        10'b0010111100:ROM_data<=18'b011111111000000000;
        10'b0010111101:ROM_data<=18'b000001100100000010;
        10'b0010111110:ROM_data<=18'b100000011111101000;
        10'b0010111111:ROM_data<=18'b111011011011111100;
        10'b0011000000:ROM_data<=18'b011111111000000000;
        10'b0011000001:ROM_data<=18'b011111110111101110;
        10'b0011000010:ROM_data<=18'b011111100111011011;
        10'b0011000011:ROM_data<=18'b011111000111001001;
        10'b0011000100:ROM_data<=18'b011111111000000000;
        10'b0011000101:ROM_data<=18'b011100011110001110;
        10'b0011000110:ROM_data<=18'b010010111100110100;
        10'b0011000111:ROM_data<=18'b000101011100000101;
        10'b0011001000:ROM_data<=18'b011111111000000000;
        10'b0011001001:ROM_data<=18'b010100110100111111;
        10'b0011001010:ROM_data<=18'b111011011100000100;
        10'b0011001011:ROM_data<=18'b100101001101111000;
        10'b0011001100:ROM_data<=18'b011111111000000000;
        10'b0011001101:ROM_data<=18'b001001111100001110;
        10'b0011001110:ROM_data<=18'b100110100101101001;
        10'b0011001111:ROM_data<=18'b100110000010010010;
        10'b0011010000:ROM_data<=18'b011111111000000000;
        10'b0011010001:ROM_data<=18'b011111011111010101;
        10'b0011010010:ROM_data<=18'b011110000110101011;
        10'b0011010011:ROM_data<=18'b011011101110000011;
        10'b0011010100:ROM_data<=18'b011111111000000000;
        10'b0011010101:ROM_data<=18'b011010111101111000;
        10'b0011010110:ROM_data<=18'b001101101100011010;
        10'b0011010111:ROM_data<=18'b111100001100000011;
        10'b0011011000:ROM_data<=18'b011111111000000000;
        10'b0011011001:ROM_data<=18'b010010010100110000;
        10'b0011011010:ROM_data<=18'b110101011100010000;
        10'b0011011011:ROM_data<=18'b100001011110111100;
        10'b0011011100:ROM_data<=18'b011111111000000000;
        10'b0011011101:ROM_data<=18'b000110111100001000;
        10'b0011011110:ROM_data<=18'b100011010110010011;
        10'b0011011111:ROM_data<=18'b101100100011001001;
        10'b0011100000:ROM_data<=18'b011111111000000000;
        10'b0011100001:ROM_data<=18'b011110101110111100;
        10'b0011100010:ROM_data<=18'b011011010101111101;
        10'b0011100011:ROM_data<=18'b010101111101001000;
        10'b0011100100:ROM_data<=18'b011111111000000000;
        10'b0011100101:ROM_data<=18'b011001001101100100;
        10'b0011100110:ROM_data<=18'b000111101100001001;
        10'b0011100111:ROM_data<=18'b110011001100010111;
        10'b0011101000:ROM_data<=18'b011111111000000000;
        10'b0011101001:ROM_data<=18'b001111101100100011;
        10'b0011101010:ROM_data<=18'b101111101100100110;
        10'b0011101011:ROM_data<=18'b100000010000000110;
        10'b0011101100:ROM_data<=18'b011111111000000000;
        10'b0011101101:ROM_data<=18'b000011111100000011;
        10'b0011101110:ROM_data<=18'b100001001111000011;
        10'b0011101111:ROM_data<=18'b110100101011101101;
        10'b0011110000:ROM_data<=18'b011111111000000000;
        10'b0011110001:ROM_data<=18'b011101101110100101;
        10'b0011110010:ROM_data<=18'b010111100101010101;
        10'b0011110011:ROM_data<=18'b001110010100011101;
        10'b0011110100:ROM_data<=18'b011111111000000000;
        10'b0011110101:ROM_data<=18'b010111000101010001;
        10'b0011110110:ROM_data<=18'b000001100100000010;
        10'b0011110111:ROM_data<=18'b101011010100111111;
        10'b0011111000:ROM_data<=18'b011111111000000000;
        10'b0011111001:ROM_data<=18'b001100111100010111;
        10'b0011111010:ROM_data<=18'b101010101101000100;
        10'b0011111011:ROM_data<=18'b100001110001001111;
        10'b0011111100:ROM_data<=18'b011111111000000000;
        10'b0011111101:ROM_data<=18'b000000110100000010;
        10'b0011111110:ROM_data<=18'b100000010111110100;
        10'b0011111111:ROM_data<=18'b111101110011111110;
        10'b0100000000:ROM_data<=18'b011111111000000000;
        10'b0100000001:ROM_data<=18'b011111110111111111;
        10'b0100000010:ROM_data<=18'b011111110111111101;
        10'b0100000011:ROM_data<=18'b011111110111111100;
        10'b0100000100:ROM_data<=18'b011111111000000000;
        10'b0100000101:ROM_data<=18'b011101010110011101;
        10'b0100000110:ROM_data<=18'b010110010101001010;
        10'b0100000111:ROM_data<=18'b001011101100010011;
        10'b0100001000:ROM_data<=18'b011111111000000000;
        10'b0100001001:ROM_data<=18'b010110011101001011;
        10'b0100001010:ROM_data<=18'b111111101100000010;
        10'b0100001011:ROM_data<=18'b101001001101010000;
        10'b0100001100:ROM_data<=18'b011111111000000000;
        10'b0100001101:ROM_data<=18'b001100000100010100;
        10'b0100001110:ROM_data<=18'b101001010101001110;
        10'b0100001111:ROM_data<=18'b100010111001100101;
        10'b0100010000:ROM_data<=18'b011111111000000000;
        10'b0100010001:ROM_data<=18'b011111101111100110;
        10'b0100010010:ROM_data<=18'b011111001111001100;
        10'b0100010011:ROM_data<=18'b011110010110110010;
        10'b0100010100:ROM_data<=18'b011111111000000000;
        10'b0100010101:ROM_data<=18'b011100000110000111;
        10'b0100010110:ROM_data<=18'b010001011100101011;
        10'b0100010111:ROM_data<=18'b000010100100000010;
        10'b0100011000:ROM_data<=18'b011111111000000000;
        10'b0100011001:ROM_data<=18'b010100000100111010;
        10'b0100011010:ROM_data<=18'b111001100100000111;
        10'b0100011011:ROM_data<=18'b100011101110001100;
        10'b0100011100:ROM_data<=18'b011111111000000000;
        10'b0100011101:ROM_data<=18'b001001000100001100;
        10'b0100011110:ROM_data<=18'b100101011101110101;
        10'b0100011111:ROM_data<=18'b100111110010100101;
        10'b0100100000:ROM_data<=18'b011111111000000000;
        10'b0100100001:ROM_data<=18'b011111001111001101;
        10'b0100100010:ROM_data<=18'b011101010110011100;
        10'b0100100011:ROM_data<=18'b011010001101101111;
        10'b0100100100:ROM_data<=18'b011111111000000000;
        10'b0100100101:ROM_data<=18'b011010011101110010;
        10'b0100100110:ROM_data<=18'b001011110100010100;
        10'b0100100111:ROM_data<=18'b111001010100000111;
        10'b0100101000:ROM_data<=18'b011111111000000000;
        10'b0100101001:ROM_data<=18'b010001100100101100;
        10'b0100101010:ROM_data<=18'b110011100100010110;
        10'b0100101011:ROM_data<=18'b100000110111010011;
        10'b0100101100:ROM_data<=18'b011111111000000000;
        10'b0100101101:ROM_data<=18'b000110000100000110;
        10'b0100101110:ROM_data<=18'b100010100110100010;
        10'b0100101111:ROM_data<=18'b101110111011010110;
        10'b0100110000:ROM_data<=18'b011111111000000000;
        10'b0100110001:ROM_data<=18'b011110011110110101;
        10'b0100110010:ROM_data<=18'b011010010101110000;
        10'b0100110011:ROM_data<=18'b010011110100111000;
        10'b0100110100:ROM_data<=18'b011111111000000000;
        10'b0100110101:ROM_data<=18'b011000100101011110;
        10'b0100110110:ROM_data<=18'b000101110100000110;
        10'b0100110111:ROM_data<=18'b110000100100100010;
        10'b0100111000:ROM_data<=18'b011111111000000000;
        10'b0100111001:ROM_data<=18'b001110110100011111;
        10'b0100111010:ROM_data<=18'b101110000100101110;
        10'b0100111011:ROM_data<=18'b100000011000011101;
        10'b0100111100:ROM_data<=18'b011111111000000000;
        10'b0100111101:ROM_data<=18'b000010111100000011;
        10'b0100111110:ROM_data<=18'b100000110111010010;
        10'b0100111111:ROM_data<=18'b110111011011110101;
        10'b0101000000:ROM_data<=18'b011111111000000000;
        10'b0101000001:ROM_data<=18'b011111110111111001;
        10'b0101000010:ROM_data<=18'b011111110111110001;
        10'b0101000011:ROM_data<=18'b011111101111101001;
        10'b0101000100:ROM_data<=18'b011111111000000000;
        10'b0101000101:ROM_data<=18'b011101000110011000;
        10'b0101000110:ROM_data<=18'b010101000101000001;
        10'b0101000111:ROM_data<=18'b001001011100001101;
        10'b0101001000:ROM_data<=18'b011111111000000000;
        10'b0101001001:ROM_data<=18'b010101110101000111;
        10'b0101001010:ROM_data<=18'b111110001100000010;
        10'b0101001011:ROM_data<=18'b100111100101011110;
        10'b0101001100:ROM_data<=18'b011111111000000000;
        10'b0101001101:ROM_data<=18'b001011010100010010;
        10'b0101001110:ROM_data<=18'b101000001101011000;
        10'b0101001111:ROM_data<=18'b100011111001110110;
        10'b0101010000:ROM_data<=18'b011111111000000000;
        10'b0101010001:ROM_data<=18'b011111100111100000;
        10'b0101010010:ROM_data<=18'b011110110111000000;
        10'b0101010011:ROM_data<=18'b011101100110100000;
        10'b0101010100:ROM_data<=18'b011111111000000000;
        10'b0101010101:ROM_data<=18'b011011101110000001;
        10'b0101010110:ROM_data<=18'b010000000100100100;
        10'b0101010111:ROM_data<=18'b000000001100000010;
        10'b0101011000:ROM_data<=18'b011111111000000000;
        10'b0101011001:ROM_data<=18'b010011011100110111;
        10'b0101011010:ROM_data<=18'b111000000100001010;
        10'b0101011011:ROM_data<=18'b100010110110011101;
        10'b0101011100:ROM_data<=18'b011111111000000000;
        10'b0101011101:ROM_data<=18'b001000010100001010;
        10'b0101011110:ROM_data<=18'b100100100110000000;
        10'b0101011111:ROM_data<=18'b101001011010110011;
        10'b0101100000:ROM_data<=18'b011111111000000000;
        10'b0101100001:ROM_data<=18'b011111000111000111;
        10'b0101100010:ROM_data<=18'b011100101110010001;
        10'b0101100011:ROM_data<=18'b011000110101100000;
        10'b0101100100:ROM_data<=18'b011111111000000000;
        10'b0101100101:ROM_data<=18'b011001111101101100;
        10'b0101100110:ROM_data<=18'b001010010100001111;
        10'b0101100111:ROM_data<=18'b110111000100001100;
        10'b0101101000:ROM_data<=18'b011111111000000000;
        10'b0101101001:ROM_data<=18'b010000111100101000;
        10'b0101101010:ROM_data<=18'b110010001100011011;
        10'b0101101011:ROM_data<=18'b100000011111100110;
        10'b0101101100:ROM_data<=18'b011111111000000000;
        10'b0101101101:ROM_data<=18'b000101010100000101;
        10'b0101101110:ROM_data<=18'b100001111110101110;
        10'b0101101111:ROM_data<=18'b110000111011100000;
        10'b0101110000:ROM_data<=18'b011111111000000000;
        10'b0101110001:ROM_data<=18'b011110001110101111;
        10'b0101110010:ROM_data<=18'b011001010101100110;
        10'b0101110011:ROM_data<=18'b010001110100101101;
        10'b0101110100:ROM_data<=18'b011111111000000000;
        10'b0101110101:ROM_data<=18'b011000000101011001;
        10'b0101110110:ROM_data<=18'b000100010100000100;
        10'b0101110111:ROM_data<=18'b101110100100101100;
        10'b0101111000:ROM_data<=18'b011111111000000000;
        10'b0101111001:ROM_data<=18'b001110001100011100;
        10'b0101111010:ROM_data<=18'b101100110100110110;
        10'b0101111011:ROM_data<=18'b100000110000110000;
        10'b0101111100:ROM_data<=18'b011111111000000000;
        10'b0101111101:ROM_data<=18'b000010001100000010;
        10'b0101111110:ROM_data<=18'b100000100111011110;
        10'b0101111111:ROM_data<=18'b111001101011111001;
        10'b0110000000:ROM_data<=18'b011111111000000000;
        10'b0110000001:ROM_data<=18'b011111110111110010;
        10'b0110000010:ROM_data<=18'b011111101111100100;
        10'b0110000011:ROM_data<=18'b011111011111010110;
        10'b0110000100:ROM_data<=18'b011111111000000000;
        10'b0110000101:ROM_data<=18'b011100101110010010;
        10'b0110000110:ROM_data<=18'b010011111100111001;
        10'b0110000111:ROM_data<=18'b000111001100001000;
        10'b0110001000:ROM_data<=18'b011111111000000000;
        10'b0110001001:ROM_data<=18'b010101010101000011;
        10'b0110001010:ROM_data<=18'b111100100100000011;
        10'b0110001011:ROM_data<=18'b100110001101101100;
        10'b0110001100:ROM_data<=18'b011111111000000000;
        10'b0110001101:ROM_data<=18'b001010100100010000;
        10'b0110001110:ROM_data<=18'b100111001101100001;
        10'b0110001111:ROM_data<=18'b100101000010000111;
        10'b0110010000:ROM_data<=18'b011111111000000000;
        10'b0110010001:ROM_data<=18'b011111100111011010;
        10'b0110010010:ROM_data<=18'b011110011110110011;
        10'b0110010011:ROM_data<=18'b011100100110001111;
        10'b0110010100:ROM_data<=18'b011111111000000000;
        10'b0110010101:ROM_data<=18'b011011001101111100;
        10'b0110010110:ROM_data<=18'b001110101100011110;
        10'b0110010111:ROM_data<=18'b111101111100000010;
        10'b0110011000:ROM_data<=18'b011111111000000000;
        10'b0110011001:ROM_data<=18'b010010110100110011;
        10'b0110011010:ROM_data<=18'b110110011100001101;
        10'b0110011011:ROM_data<=18'b100001111110101111;
        10'b0110011100:ROM_data<=18'b011111111000000000;
        10'b0110011101:ROM_data<=18'b000111100100001001;
        10'b0110011110:ROM_data<=18'b100011110110001011;
        10'b0110011111:ROM_data<=18'b101011001011000000;
        10'b0110100000:ROM_data<=18'b011111111000000000;
        10'b0110100001:ROM_data<=18'b011110110111000001;
        10'b0110100010:ROM_data<=18'b011011111110000110;
        10'b0110100011:ROM_data<=18'b010111001101010010;
        10'b0110100100:ROM_data<=18'b011111111000000000;
        10'b0110100101:ROM_data<=18'b011001011101100111;
        10'b0110100110:ROM_data<=18'b001000111100001100;
        10'b0110100111:ROM_data<=18'b110100110100010010;
        10'b0110101000:ROM_data<=18'b011111111000000000;
        10'b0110101001:ROM_data<=18'b010000001100100101;
        10'b0110101010:ROM_data<=18'b110000110100100001;
        10'b0110101011:ROM_data<=18'b100000010111111001;
        10'b0110101100:ROM_data<=18'b011111111000000000;
        10'b0110101101:ROM_data<=18'b000100011100000100;
        10'b0110101110:ROM_data<=18'b100001100110111001;
        10'b0110101111:ROM_data<=18'b110011000011101000;
        10'b0110110000:ROM_data<=18'b011111111000000000;
        10'b0110110001:ROM_data<=18'b011101111110101001;
        10'b0110110010:ROM_data<=18'b011000011101011100;
        10'b0110110011:ROM_data<=18'b001111111100100011;
        10'b0110110100:ROM_data<=18'b011111111000000000;
        10'b0110110101:ROM_data<=18'b010111011101010100;
        10'b0110110110:ROM_data<=18'b000010101100000010;
        10'b0110110111:ROM_data<=18'b101100101100110111;
        10'b0110111000:ROM_data<=18'b011111111000000000;
        10'b0110111001:ROM_data<=18'b001101011100011001;
        10'b0110111010:ROM_data<=18'b101011100100111101;
        10'b0110111011:ROM_data<=18'b100001010001000010;
        10'b0110111100:ROM_data<=18'b011111111000000000;
        10'b0110111101:ROM_data<=18'b000001010100000010;
        10'b0110111110:ROM_data<=18'b100000010111101011;
        10'b0110111111:ROM_data<=18'b111100000011111100;
        10'b0111000000:ROM_data<=18'b011111111000000000;
        10'b0111000001:ROM_data<=18'b011111110111101100;
        10'b0111000010:ROM_data<=18'b011111011111011000;
        10'b0111000011:ROM_data<=18'b011110111111000100;
        10'b0111000100:ROM_data<=18'b011111111000000000;
        10'b0111000101:ROM_data<=18'b011100011110001100;
        10'b0111000110:ROM_data<=18'b010010101100110010;
        10'b0111000111:ROM_data<=18'b000100110100000100;
        10'b0111001000:ROM_data<=18'b011111111000000000;
        10'b0111001001:ROM_data<=18'b010100101100111110;
        10'b0111001010:ROM_data<=18'b111011000100000101;
        10'b0111001011:ROM_data<=18'b100100111101111100;
        10'b0111001100:ROM_data<=18'b011111111000000000;
        10'b0111001101:ROM_data<=18'b001001110100001110;
        10'b0111001110:ROM_data<=18'b100110010101101011;
        10'b0111001111:ROM_data<=18'b100110011010010110;
        10'b0111010000:ROM_data<=18'b011111111000000000;
        10'b0111010001:ROM_data<=18'b011111010111010011;
        10'b0111010010:ROM_data<=18'b011101111110101000;
        10'b0111010011:ROM_data<=18'b011011011101111111;
        10'b0111010100:ROM_data<=18'b011111111000000000;
        10'b0111010101:ROM_data<=18'b011010110101110111;
        10'b0111010110:ROM_data<=18'b001101010100011001;
        10'b0111010111:ROM_data<=18'b111011101100000100;
        10'b0111011000:ROM_data<=18'b011111111000000000;
        10'b0111011001:ROM_data<=18'b010010001100101111;
        10'b0111011010:ROM_data<=18'b110101000100010001;
        10'b0111011011:ROM_data<=18'b100001010111000001;
        10'b0111011100:ROM_data<=18'b011111111000000000;
        10'b0111011101:ROM_data<=18'b000110110100000111;
        10'b0111011110:ROM_data<=18'b100011001110010110;
        10'b0111011111:ROM_data<=18'b101100111011001011;
        10'b0111100000:ROM_data<=18'b011111111000000000;
        10'b0111100001:ROM_data<=18'b011110101110111011;
        10'b0111100010:ROM_data<=18'b011011001101111011;
        10'b0111100011:ROM_data<=18'b010101100101000101;
        10'b0111100100:ROM_data<=18'b011111111000000000;
        10'b0111100101:ROM_data<=18'b011001000101100010;
        10'b0111100110:ROM_data<=18'b000111010100001000;
        10'b0111100111:ROM_data<=18'b110010101100011001;
        10'b0111101000:ROM_data<=18'b011111111000000000;
        10'b0111101001:ROM_data<=18'b001111100100100010;
        10'b0111101010:ROM_data<=18'b101111011100100111;
        10'b0111101011:ROM_data<=18'b100000010000001010;
        10'b0111101100:ROM_data<=18'b011111111000000000;
        10'b0111101101:ROM_data<=18'b000011101100000011;
        10'b0111101110:ROM_data<=18'b100001000111000110;
        10'b0111101111:ROM_data<=18'b110101001011101111;
        10'b0111110000:ROM_data<=18'b011111111000000000;
        10'b0111110001:ROM_data<=18'b011101101110100011;
        10'b0111110010:ROM_data<=18'b010111010101010011;
        10'b0111110011:ROM_data<=18'b001101110100011011;
        10'b0111110100:ROM_data<=18'b011111111000000000;
        10'b0111110101:ROM_data<=18'b010110111101010000;
        10'b0111110110:ROM_data<=18'b000001001100000010;
        10'b0111110111:ROM_data<=18'b101010110101000011;
        10'b0111111000:ROM_data<=18'b011111111000000000;
        10'b0111111001:ROM_data<=18'b001100101100010111;
        10'b0111111010:ROM_data<=18'b101010011101000110;
        10'b0111111011:ROM_data<=18'b100010000001010100;
        10'b0111111100:ROM_data<=18'b011111111000000000;
        10'b0111111101:ROM_data<=18'b000000100100000010;
        10'b0111111110:ROM_data<=18'b100000010111110111;
        10'b0111111111:ROM_data<=18'b111110010011111110;
        10'b1000000000:ROM_data<=18'b011111111000000000;
        10'b1000000001:ROM_data<=18'b011111110111111101;
        10'b1000000010:ROM_data<=18'b011111110111111010;
        10'b1000000011:ROM_data<=18'b011111110111110111;
        10'b1000000100:ROM_data<=18'b011111111000000000;
        10'b1000000101:ROM_data<=18'b011101010110011100;
        10'b1000000110:ROM_data<=18'b010101111101001000;
        10'b1000000111:ROM_data<=18'b001011000100010001;
        10'b1000001000:ROM_data<=18'b011111111000000000;
        10'b1000001001:ROM_data<=18'b010110010101001010;
        10'b1000001010:ROM_data<=18'b111111010100000010;
        10'b1000001011:ROM_data<=18'b101000110101010011;
        10'b1000001100:ROM_data<=18'b011111111000000000;
        10'b1000001101:ROM_data<=18'b001011110100010100;
        10'b1000001110:ROM_data<=18'b101001000101010001;
        10'b1000001111:ROM_data<=18'b100011001001101010;
        10'b1000010000:ROM_data<=18'b011111111000000000;
        10'b1000010001:ROM_data<=18'b011111101111100100;
        10'b1000010010:ROM_data<=18'b011111000111001001;
        10'b1000010011:ROM_data<=18'b011110001110101110;
        10'b1000010100:ROM_data<=18'b011111111000000000;
        10'b1000010101:ROM_data<=18'b011011111110000110;
        10'b1000010110:ROM_data<=18'b010001000100101001;
        10'b1000010111:ROM_data<=18'b000001111100000010;
        10'b1000011000:ROM_data<=18'b011111111000000000;
        10'b1000011001:ROM_data<=18'b010011111100111001;
        10'b1000011010:ROM_data<=18'b111001001100001000;
        10'b1000011011:ROM_data<=18'b100011011110010001;
        10'b1000011100:ROM_data<=18'b011111111000000000;
        10'b1000011101:ROM_data<=18'b001000111100001100;
        10'b1000011110:ROM_data<=18'b100101001101111000;
        10'b1000011111:ROM_data<=18'b101000001010101000;
        10'b1000100000:ROM_data<=18'b011111111000000000;
        10'b1000100001:ROM_data<=18'b011111001111001100;
        10'b1000100010:ROM_data<=18'b011101001110011001;
        10'b1000100011:ROM_data<=18'b011001110101101011;
        10'b1000100100:ROM_data<=18'b011111111000000000;
        10'b1000100101:ROM_data<=18'b011010010101110000;
        10'b1000100110:ROM_data<=18'b001011011100010011;
        10'b1000100111:ROM_data<=18'b111000110100001000;
        10'b1000101000:ROM_data<=18'b011111111000000000;
        10'b1000101001:ROM_data<=18'b010001011100101011;
        10'b1000101010:ROM_data<=18'b110011001100010111;
        10'b1000101011:ROM_data<=18'b100000101111011000;
        10'b1000101100:ROM_data<=18'b011111111000000000;
        10'b1000101101:ROM_data<=18'b000101110100000110;
        10'b1000101110:ROM_data<=18'b100010011110100101;
        10'b1000101111:ROM_data<=18'b101111011011011001;
        10'b1000110000:ROM_data<=18'b011111111000000000;
        10'b1000110001:ROM_data<=18'b011110011110110011;
        10'b1000110010:ROM_data<=18'b011010000101101110;
        10'b1000110011:ROM_data<=18'b010011010100110110;
        10'b1000110100:ROM_data<=18'b011111111000000000;
        10'b1000110101:ROM_data<=18'b011000011101011100;
        10'b1000110110:ROM_data<=18'b000101011100000101;
        10'b1000110111:ROM_data<=18'b110000000100100100;
        10'b1000111000:ROM_data<=18'b011111111000000000;
        10'b1000111001:ROM_data<=18'b001110101100011110;
        10'b1000111010:ROM_data<=18'b101101110100110000;
        10'b1000111011:ROM_data<=18'b100000100000100010;
        10'b1000111100:ROM_data<=18'b011111111000000000;
        10'b1000111101:ROM_data<=18'b000010101100000010;
        10'b1000111110:ROM_data<=18'b100000101111010101;
        10'b1000111111:ROM_data<=18'b111000000011110110;
        10'b1001000000:ROM_data<=18'b011111111000000000;
        10'b1001000001:ROM_data<=18'b011111110111110111;
        10'b1001000010:ROM_data<=18'b011111110111101110;
        10'b1001000011:ROM_data<=18'b011111101111100100;
        10'b1001000100:ROM_data<=18'b011111111000000000;
        10'b1001000101:ROM_data<=18'b011100111110010110;
        10'b1001000110:ROM_data<=18'b010100110100111111;
        10'b1001000111:ROM_data<=18'b001000111100001100;
        10'b1001001000:ROM_data<=18'b011111111000000000;
        10'b1001001001:ROM_data<=18'b010101101101000110;
        10'b1001001010:ROM_data<=18'b111101110100000010;
        10'b1001001011:ROM_data<=18'b100111001101100001;
        10'b1001001100:ROM_data<=18'b011111111000000000;
        10'b1001001101:ROM_data<=18'b001011000100010001;
        10'b1001001110:ROM_data<=18'b100111111101011010;
        10'b1001001111:ROM_data<=18'b100100001001111010;
        10'b1001010000:ROM_data<=18'b011111111000000000;
        10'b1001010001:ROM_data<=18'b011111100111011110;
        10'b1001010010:ROM_data<=18'b011110101110111100;
        10'b1001010011:ROM_data<=18'b011101010110011100;
        10'b1001010100:ROM_data<=18'b011111111000000000;
        10'b1001010101:ROM_data<=18'b011011100110000000;
        10'b1001010110:ROM_data<=18'b001111101100100011;
        10'b1001010111:ROM_data<=18'b111111101100000010;
        10'b1001011000:ROM_data<=18'b011111111000000000;
        10'b1001011001:ROM_data<=18'b010011010100110110;
        10'b1001011010:ROM_data<=18'b110111100100001011;
        10'b1001011011:ROM_data<=18'b100010100110100010;
        10'b1001011100:ROM_data<=18'b011111111000000000;
        10'b1001011101:ROM_data<=18'b001000000100001010;
        10'b1001011110:ROM_data<=18'b100100011110000011;
        10'b1001011111:ROM_data<=18'b101001110010110110;
        10'b1001100000:ROM_data<=18'b011111111000000000;
        10'b1001100001:ROM_data<=18'b011111000111000110;
        10'b1001100010:ROM_data<=18'b011100011110001110;
        10'b1001100011:ROM_data<=18'b011000011101011100;
        10'b1001100100:ROM_data<=18'b011111111000000000;
        10'b1001100101:ROM_data<=18'b011001110101101011;
        10'b1001100110:ROM_data<=18'b001001111100001110;
        10'b1001100111:ROM_data<=18'b110110011100001101;
        10'b1001101000:ROM_data<=18'b011111111000000000;
        10'b1001101001:ROM_data<=18'b010000101100100111;
        10'b1001101010:ROM_data<=18'b110001110100011101;
        10'b1001101011:ROM_data<=18'b100000010111101011;
        10'b1001101100:ROM_data<=18'b011111111000000000;
        10'b1001101101:ROM_data<=18'b000101000100000101;
        10'b1001101110:ROM_data<=18'b100001110110110001;
        10'b1001101111:ROM_data<=18'b110001011011100010;
        10'b1001110000:ROM_data<=18'b011111111000000000;
        10'b1001110001:ROM_data<=18'b011110001110101110;
        10'b1001110010:ROM_data<=18'b011001001101100100;
        10'b1001110011:ROM_data<=18'b010001011100101011;
        10'b1001110100:ROM_data<=18'b011111111000000000;
        10'b1001110101:ROM_data<=18'b010111111101011000;
        10'b1001110110:ROM_data<=18'b000011111100000011;
        10'b1001110111:ROM_data<=18'b101110000100101110;
        10'b1001111000:ROM_data<=18'b011111111000000000;
        10'b1001111001:ROM_data<=18'b001101111100011011;
        10'b1001111010:ROM_data<=18'b101100100100110111;
        10'b1001111011:ROM_data<=18'b100000111000110100;
        10'b1001111100:ROM_data<=18'b011111111000000000;
        10'b1001111101:ROM_data<=18'b000001111100000010;
        10'b1001111110:ROM_data<=18'b100000011111100001;
        10'b1001111111:ROM_data<=18'b111010010011111010;
        10'b1010000000:ROM_data<=18'b011111111000000000;
        10'b1010000001:ROM_data<=18'b011111110111110001;
        10'b1010000010:ROM_data<=18'b011111101111100001;
        10'b1010000011:ROM_data<=18'b011111010111010010;
        10'b1010000100:ROM_data<=18'b011111111000000000;
        10'b1010000101:ROM_data<=18'b011100101110010001;
        10'b1010000110:ROM_data<=18'b010011100100110111;
        10'b1010000111:ROM_data<=18'b000110100100000111;
        10'b1010001000:ROM_data<=18'b011111111000000000;
        10'b1010001001:ROM_data<=18'b010101000101000001;
        10'b1010001010:ROM_data<=18'b111100001100000011;
        10'b1010001011:ROM_data<=18'b100101110101110000;
        10'b1010001100:ROM_data<=18'b011111111000000000;
        10'b1010001101:ROM_data<=18'b001010010100001111;
        10'b1010001110:ROM_data<=18'b100110111101100100;
        10'b1010001111:ROM_data<=18'b100101011010001011;
        10'b1010010000:ROM_data<=18'b011111111000000000;
        10'b1010010001:ROM_data<=18'b011111011111011000;
        10'b1010010010:ROM_data<=18'b011110010110110001;
        10'b1010010011:ROM_data<=18'b011100010110001011;
        10'b1010010100:ROM_data<=18'b011111111000000000;
        10'b1010010101:ROM_data<=18'b011011001101111011;
        10'b1010010110:ROM_data<=18'b001110010100011101;
        10'b1010010111:ROM_data<=18'b111101011100000010;
        10'b1010011000:ROM_data<=18'b011111111000000000;
        10'b1010011001:ROM_data<=18'b010010101100110010;
        10'b1010011010:ROM_data<=18'b110110001100001110;
        10'b1010011011:ROM_data<=18'b100001101110110011;
        10'b1010011100:ROM_data<=18'b011111111000000000;
        10'b1010011101:ROM_data<=18'b000111010100001000;
        10'b1010011110:ROM_data<=18'b100011101110001110;
        10'b1010011111:ROM_data<=18'b101011100011000011;
        10'b1010100000:ROM_data<=18'b011111111000000000;
        10'b1010100001:ROM_data<=18'b011110110111000000;
        10'b1010100010:ROM_data<=18'b011011101110000011;
        10'b1010100011:ROM_data<=18'b010110110101001110;
        10'b1010100100:ROM_data<=18'b011111111000000000;
        10'b1010100101:ROM_data<=18'b011001010101100110;
        10'b1010100110:ROM_data<=18'b001000100100001011;
        10'b1010100111:ROM_data<=18'b110100010100010100;
        10'b1010101000:ROM_data<=18'b011111111000000000;
        10'b1010101001:ROM_data<=18'b010000000100100100;
        10'b1010101010:ROM_data<=18'b110000011100100011;
        10'b1010101011:ROM_data<=18'b100000010111111101;
        10'b1010101100:ROM_data<=18'b011111111000000000;
        10'b1010101101:ROM_data<=18'b000100010100000100;
        10'b1010101110:ROM_data<=18'b100001011110111100;
        10'b1010101111:ROM_data<=18'b110011100011101010;
        10'b1010110000:ROM_data<=18'b011111111000000000;
        10'b1010110001:ROM_data<=18'b011101111110101000;
        10'b1010110010:ROM_data<=18'b011000001101011010;
        10'b1010110011:ROM_data<=18'b001111010100100001;
        10'b1010110100:ROM_data<=18'b011111111000000000;
        10'b1010110101:ROM_data<=18'b010111010101010011;
        10'b1010110110:ROM_data<=18'b000010010100000010;
        10'b1010110111:ROM_data<=18'b101100001100111001;
        10'b1010111000:ROM_data<=18'b011111111000000000;
        10'b1010111001:ROM_data<=18'b001101010100011001;
        10'b1010111010:ROM_data<=18'b101011010100111111;
        10'b1010111011:ROM_data<=18'b100001100001000111;
        10'b1010111100:ROM_data<=18'b011111111000000000;
        10'b1010111101:ROM_data<=18'b000001001100000010;
        10'b1010111110:ROM_data<=18'b100000010111101110;
        10'b1010111111:ROM_data<=18'b111100100011111101;
        10'b1011000000:ROM_data<=18'b011111111000000000;
        10'b1011000001:ROM_data<=18'b011111110111101011;
        10'b1011000010:ROM_data<=18'b011111011111010101;
        10'b1011000011:ROM_data<=18'b011110110111000000;
        10'b1011000100:ROM_data<=18'b011111111000000000;
        10'b1011000101:ROM_data<=18'b011100010110001011;
        10'b1011000110:ROM_data<=18'b010010010100110000;
        10'b1011000111:ROM_data<=18'b000100010100000100;
        10'b1011001000:ROM_data<=18'b011111111000000000;
        10'b1011001001:ROM_data<=18'b010100100100111101;
        10'b1011001010:ROM_data<=18'b111010101100000101;
        10'b1011001011:ROM_data<=18'b100100100110000000;
        10'b1011001100:ROM_data<=18'b011111111000000000;
        10'b1011001101:ROM_data<=18'b001001101100001101;
        10'b1011001110:ROM_data<=18'b100110000101101110;
        10'b1011001111:ROM_data<=18'b100110110010011010;
        10'b1011010000:ROM_data<=18'b011111111000000000;
        10'b1011010001:ROM_data<=18'b011111010111010010;
        10'b1011010010:ROM_data<=18'b011101101110100101;
        10'b1011010011:ROM_data<=18'b011011001101111011;
        10'b1011010100:ROM_data<=18'b011111111000000000;
        10'b1011010101:ROM_data<=18'b011010101101110101;
        10'b1011010110:ROM_data<=18'b001100111100010111;
        10'b1011010111:ROM_data<=18'b111011000100000101;
        10'b1011011000:ROM_data<=18'b011111111000000000;
        10'b1011011001:ROM_data<=18'b010010000100101110;
        10'b1011011010:ROM_data<=18'b110100101100010011;
        10'b1011011011:ROM_data<=18'b100001000111000110;
        10'b1011011100:ROM_data<=18'b011111111000000000;
        10'b1011011101:ROM_data<=18'b000110100100000111;
        10'b1011011110:ROM_data<=18'b100010111110011001;
        10'b1011011111:ROM_data<=18'b101101011011001110;
        10'b1011100000:ROM_data<=18'b011111111000000000;
        10'b1011100001:ROM_data<=18'b011110100110111001;
        10'b1011100010:ROM_data<=18'b011010111101111000;
        10'b1011100011:ROM_data<=18'b010101000101000001;
        10'b1011100100:ROM_data<=18'b011111111000000000;
        10'b1011100101:ROM_data<=18'b011000111101100001;
        10'b1011100110:ROM_data<=18'b000110111100001000;
        10'b1011100111:ROM_data<=18'b110010001100011011;
        10'b1011101000:ROM_data<=18'b011111111000000000;
        10'b1011101001:ROM_data<=18'b001111010100100001;
        10'b1011101010:ROM_data<=18'b101111000100101001;
        10'b1011101011:ROM_data<=18'b100000010000001111;
        10'b1011101100:ROM_data<=18'b011111111000000000;
        10'b1011101101:ROM_data<=18'b000011100100000011;
        10'b1011101110:ROM_data<=18'b100001000111001001;
        10'b1011101111:ROM_data<=18'b110101110011110001;
        10'b1011110000:ROM_data<=18'b011111111000000000;
        10'b1011110001:ROM_data<=18'b011101100110100010;
        10'b1011110010:ROM_data<=18'b010111000101010001;
        10'b1011110011:ROM_data<=18'b001101010100011001;
        10'b1011110100:ROM_data<=18'b011111111000000000;
        10'b1011110101:ROM_data<=18'b010110110101001110;
        10'b1011110110:ROM_data<=18'b000000110100000010;
        10'b1011110111:ROM_data<=18'b101010011101000110;
        10'b1011111000:ROM_data<=18'b011111111000000000;
        10'b1011111001:ROM_data<=18'b001100100100010110;
        10'b1011111010:ROM_data<=18'b101010001101001000;
        10'b1011111011:ROM_data<=18'b100010001001011000;
        10'b1011111100:ROM_data<=18'b011111111000000000;
        10'b1011111101:ROM_data<=18'b000000011100000010;
        10'b1011111110:ROM_data<=18'b100000010111111010;
        10'b1011111111:ROM_data<=18'b111110111011111110;
        10'b1100000000:ROM_data<=18'b011111111000000000;
        10'b1100000001:ROM_data<=18'b011111110111111100;
        10'b1100000010:ROM_data<=18'b011111110111110111;
        10'b1100000011:ROM_data<=18'b011111110111110010;
        10'b1100000100:ROM_data<=18'b011111111000000000;
        10'b1100000101:ROM_data<=18'b011101001110011011;
        10'b1100000110:ROM_data<=18'b010101101101000110;
        10'b1100000111:ROM_data<=18'b001010100100010000;
        10'b1100001000:ROM_data<=18'b011111111000000000;
        10'b1100001001:ROM_data<=18'b010110000101001001;
        10'b1100001010:ROM_data<=18'b111110111100000010;
        10'b1100001011:ROM_data<=18'b101000011101010110;
        10'b1100001100:ROM_data<=18'b011111111000000000;
        10'b1100001101:ROM_data<=18'b001011101100010011;
        10'b1100001110:ROM_data<=18'b101000110101010011;
        10'b1100001111:ROM_data<=18'b100011011001101110;
        10'b1100010000:ROM_data<=18'b011111111000000000;
        10'b1100010001:ROM_data<=18'b011111101111100011;
        10'b1100010010:ROM_data<=18'b011111000111000110;
        10'b1100010011:ROM_data<=18'b011101111110101001;
        10'b1100010100:ROM_data<=18'b011111111000000000;
        10'b1100010101:ROM_data<=18'b011011110110000100;
        10'b1100010110:ROM_data<=18'b010000101100100111;
        10'b1100010111:ROM_data<=18'b000001010100000010;
        10'b1100011000:ROM_data<=18'b011111111000000000;
        10'b1100011001:ROM_data<=18'b010011110100111000;
        10'b1100011010:ROM_data<=18'b111000110100001000;
        10'b1100011011:ROM_data<=18'b100011001110010101;
        10'b1100011100:ROM_data<=18'b011111111000000000;
        10'b1100011101:ROM_data<=18'b001000101100001011;
        10'b1100011110:ROM_data<=18'b100100111101111011;
        10'b1100011111:ROM_data<=18'b101000101010101100;
        10'b1100100000:ROM_data<=18'b011111111000000000;
        10'b1100100001:ROM_data<=18'b011111001111001010;
        10'b1100100010:ROM_data<=18'b011100111110010110;
        10'b1100100011:ROM_data<=18'b011001011101100111;
        10'b1100100100:ROM_data<=18'b011111111000000000;
        10'b1100100101:ROM_data<=18'b011010001101101111;
        10'b1100100110:ROM_data<=18'b001011000100010001;
        10'b1100100111:ROM_data<=18'b111000001100001010;
        10'b1100101000:ROM_data<=18'b011111111000000000;
        10'b1100101001:ROM_data<=18'b010001001100101010;
        10'b1100101010:ROM_data<=18'b110010110100011001;
        10'b1100101011:ROM_data<=18'b100000100111011101;
        10'b1100101100:ROM_data<=18'b011111111000000000;
        10'b1100101101:ROM_data<=18'b000101101100000110;
        10'b1100101110:ROM_data<=18'b100010001110101000;
        10'b1100101111:ROM_data<=18'b101111111011011011;
        10'b1100110000:ROM_data<=18'b011111111000000000;
        10'b1100110001:ROM_data<=18'b011110010110110010;
        10'b1100110010:ROM_data<=18'b011001110101101011;
        10'b1100110011:ROM_data<=18'b010010110100110011;
        10'b1100110100:ROM_data<=18'b011111111000000000;
        10'b1100110101:ROM_data<=18'b011000010101011011;
        10'b1100110110:ROM_data<=18'b000101000100000101;
        10'b1100110111:ROM_data<=18'b101111100100100111;
        10'b1100111000:ROM_data<=18'b011111111000000000;
        10'b1100111001:ROM_data<=18'b001110100100011101;
        10'b1100111010:ROM_data<=18'b101101011100110010;
        10'b1100111011:ROM_data<=18'b100000100000100110;
        10'b1100111100:ROM_data<=18'b011111111000000000;
        10'b1100111101:ROM_data<=18'b000010100100000010;
        10'b1100111110:ROM_data<=18'b100000101111011000;
        10'b1100111111:ROM_data<=18'b111000100011110111;
        10'b1101000000:ROM_data<=18'b011111111000000000;
        10'b1101000001:ROM_data<=18'b011111110111110110;
        10'b1101000010:ROM_data<=18'b011111110111101011;
        10'b1101000011:ROM_data<=18'b011111100111100000;
        10'b1101000100:ROM_data<=18'b011111111000000000;
        10'b1101000101:ROM_data<=18'b011100111110010101;
        10'b1101000110:ROM_data<=18'b010100100100111101;
        10'b1101000111:ROM_data<=18'b001000010100001010;
        10'b1101001000:ROM_data<=18'b011111111000000000;
        10'b1101001001:ROM_data<=18'b010101100101000101;
        10'b1101001010:ROM_data<=18'b111101011100000010;
        10'b1101001011:ROM_data<=18'b100110111101100101;
        10'b1101001100:ROM_data<=18'b011111111000000000;
        10'b1101001101:ROM_data<=18'b001010111100010001;
        10'b1101001110:ROM_data<=18'b100111101101011100;
        10'b1101001111:ROM_data<=18'b100100011001111111;
        10'b1101010000:ROM_data<=18'b011111111000000000;
        10'b1101010001:ROM_data<=18'b011111100111011101;
        10'b1101010010:ROM_data<=18'b011110100110111001;
        10'b1101010011:ROM_data<=18'b011101000110011000;
        10'b1101010100:ROM_data<=18'b011111111000000000;
        10'b1101010101:ROM_data<=18'b011011011101111111;
        10'b1101010110:ROM_data<=18'b001111010100100001;
        10'b1101010111:ROM_data<=18'b111111001100000010;
        10'b1101011000:ROM_data<=18'b011111111000000000;
        10'b1101011001:ROM_data<=18'b010011001100110101;
        10'b1101011010:ROM_data<=18'b110111001100001100;
        10'b1101011011:ROM_data<=18'b100010010110100110;
        10'b1101011100:ROM_data<=18'b011111111000000000;
        10'b1101011101:ROM_data<=18'b000111111100001010;
        10'b1101011110:ROM_data<=18'b100100001110000110;
        10'b1101011111:ROM_data<=18'b101010010010111001;
        10'b1101100000:ROM_data<=18'b011111111000000000;
        10'b1101100001:ROM_data<=18'b011110111111000100;
        10'b1101100010:ROM_data<=18'b011100010110001011;
        10'b1101100011:ROM_data<=18'b011000000101011001;
        10'b1101100100:ROM_data<=18'b011111111000000000;
        10'b1101100101:ROM_data<=18'b011001101101101010;
        10'b1101100110:ROM_data<=18'b001001101100001101;
        10'b1101100111:ROM_data<=18'b110101111100001111;
        10'b1101101000:ROM_data<=18'b011111111000000000;
        10'b1101101001:ROM_data<=18'b010000100100100111;
        10'b1101101010:ROM_data<=18'b110001011100011110;
        10'b1101101011:ROM_data<=18'b100000010111101111;
        10'b1101101100:ROM_data<=18'b011111111000000000;
        10'b1101101101:ROM_data<=18'b000100110100000100;
        10'b1101101110:ROM_data<=18'b100001101110110011;
        10'b1101101111:ROM_data<=18'b110001111011100100;
        10'b1101110000:ROM_data<=18'b011111111000000000;
        10'b1101110001:ROM_data<=18'b011110000110101100;
        10'b1101110010:ROM_data<=18'b011000111101100001;
        10'b1101110011:ROM_data<=18'b010000111100101000;
        10'b1101110100:ROM_data<=18'b011111111000000000;
        10'b1101110101:ROM_data<=18'b010111101101010110;
        10'b1101110110:ROM_data<=18'b000011100100000011;
        10'b1101110111:ROM_data<=18'b101101100100110001;
        10'b1101111000:ROM_data<=18'b011111111000000000;
        10'b1101111001:ROM_data<=18'b001101110100011011;
        10'b1101111010:ROM_data<=18'b101100001100111001;
        10'b1101111011:ROM_data<=18'b100001000000111001;
        10'b1101111100:ROM_data<=18'b011111111000000000;
        10'b1101111101:ROM_data<=18'b000001110100000010;
        10'b1101111110:ROM_data<=18'b100000011111100100;
        10'b1101111111:ROM_data<=18'b111010110011111011;
        10'b1110000000:ROM_data<=18'b011111111000000000;
        10'b1110000001:ROM_data<=18'b011111110111101111;
        10'b1110000010:ROM_data<=18'b011111100111011110;
        10'b1110000011:ROM_data<=18'b011111001111001101;
        10'b1110000100:ROM_data<=18'b011111111000000000;
        10'b1110000101:ROM_data<=18'b011100100110001111;
        10'b1110000110:ROM_data<=18'b010011010100110110;
        10'b1110000111:ROM_data<=18'b000110000100000110;
        10'b1110001000:ROM_data<=18'b011111111000000000;
        10'b1110001001:ROM_data<=18'b010100111101000000;
        10'b1110001010:ROM_data<=18'b111011110100000100;
        10'b1110001011:ROM_data<=18'b100101100101110100;
        10'b1110001100:ROM_data<=18'b011111111000000000;
        10'b1110001101:ROM_data<=18'b001010001100001111;
        10'b1110001110:ROM_data<=18'b100110110101100110;
        10'b1110001111:ROM_data<=18'b100101101010001110;
        10'b1110010000:ROM_data<=18'b011111111000000000;
        10'b1110010001:ROM_data<=18'b011111011111010110;
        10'b1110010010:ROM_data<=18'b011110001110101110;
        10'b1110010011:ROM_data<=18'b011100000110000111;
        10'b1110010100:ROM_data<=18'b011111111000000000;
        10'b1110010101:ROM_data<=18'b011011000101111001;
        10'b1110010110:ROM_data<=18'b001101111100011011;
        10'b1110010111:ROM_data<=18'b111100110100000011;
        10'b1110011000:ROM_data<=18'b011111111000000000;
        10'b1110011001:ROM_data<=18'b010010100100110001;
        10'b1110011010:ROM_data<=18'b110101110100001111;
        10'b1110011011:ROM_data<=18'b100001100110111000;
        10'b1110011100:ROM_data<=18'b011111111000000000;
        10'b1110011101:ROM_data<=18'b000111001100001000;
        10'b1110011110:ROM_data<=18'b100011011110010001;
        10'b1110011111:ROM_data<=18'b101100000011000110;
        10'b1110100000:ROM_data<=18'b011111111000000000;
        10'b1110100001:ROM_data<=18'b011110110110111110;
        10'b1110100010:ROM_data<=18'b011011100110000000;
        10'b1110100011:ROM_data<=18'b010110011101001011;
        10'b1110100100:ROM_data<=18'b011111111000000000;
        10'b1110100101:ROM_data<=18'b011001001101100101;
        10'b1110100110:ROM_data<=18'b001000000100001010;
        10'b1110100111:ROM_data<=18'b110011101100010110;
        10'b1110101000:ROM_data<=18'b011111111000000000;
        10'b1110101001:ROM_data<=18'b001111111100100011;
        10'b1110101010:ROM_data<=18'b110000000100100100;
        10'b1110101011:ROM_data<=18'b100000010000000001;
        10'b1110101100:ROM_data<=18'b011111111000000000;
        10'b1110101101:ROM_data<=18'b000100000100000100;
        10'b1110101110:ROM_data<=18'b100001010111000000;
        10'b1110101111:ROM_data<=18'b110100000011101100;
        10'b1110110000:ROM_data<=18'b011111111000000000;
        10'b1110110001:ROM_data<=18'b011101110110100110;
        10'b1110110010:ROM_data<=18'b010111111101011000;
        10'b1110110011:ROM_data<=18'b001110110100011111;
        10'b1110110100:ROM_data<=18'b011111111000000000;
        10'b1110110101:ROM_data<=18'b010111001101010010;
        10'b1110110110:ROM_data<=18'b000001111100000010;
        10'b1110110111:ROM_data<=18'b101011110100111100;
        10'b1110111000:ROM_data<=18'b011111111000000000;
        10'b1110111001:ROM_data<=18'b001101000100011000;
        10'b1110111010:ROM_data<=18'b101011000101000001;
        10'b1110111011:ROM_data<=18'b100001101001001011;
        10'b1110111100:ROM_data<=18'b011111111000000000;
        10'b1110111101:ROM_data<=18'b000000111100000010;
        10'b1110111110:ROM_data<=18'b100000010111110001;
        10'b1110111111:ROM_data<=18'b111101001011111101;
        10'b1111000000:ROM_data<=18'b011111111000000000;
        10'b1111000001:ROM_data<=18'b011111101111101001;
        10'b1111000010:ROM_data<=18'b011111010111010010;
        10'b1111000011:ROM_data<=18'b011110101110111011;
        10'b1111000100:ROM_data<=18'b011111111000000000;
        10'b1111000101:ROM_data<=18'b011100001110001010;
        10'b1111000110:ROM_data<=18'b010010000100101110;
        10'b1111000111:ROM_data<=18'b000011101100000011;
        10'b1111001000:ROM_data<=18'b011111111000000000;
        10'b1111001001:ROM_data<=18'b010100010100111100;
        10'b1111001010:ROM_data<=18'b111010010100000110;
        10'b1111001011:ROM_data<=18'b100100010110000100;
        10'b1111001100:ROM_data<=18'b011111111000000000;
        10'b1111001101:ROM_data<=18'b001001011100001101;
        10'b1111001110:ROM_data<=18'b100101110101110000;
        10'b1111001111:ROM_data<=18'b100111000010011110;
        10'b1111010000:ROM_data<=18'b011111111000000000;
        10'b1111010001:ROM_data<=18'b011111010111010000;
        10'b1111010010:ROM_data<=18'b011101100110100010;
        10'b1111010011:ROM_data<=18'b011010110101110111;
        10'b1111010100:ROM_data<=18'b011111111000000000;
        10'b1111010101:ROM_data<=18'b011010100101110100;
        10'b1111010110:ROM_data<=18'b001100100100010110;
        10'b1111010111:ROM_data<=18'b111010011100000110;
        10'b1111011000:ROM_data<=18'b011111111000000000;
        10'b1111011001:ROM_data<=18'b010001110100101101;
        10'b1111011010:ROM_data<=18'b110100010100010100;
        10'b1111011011:ROM_data<=18'b100000111111001010;
        10'b1111011100:ROM_data<=18'b011111111000000000;
        10'b1111011101:ROM_data<=18'b000110011100000111;
        10'b1111011110:ROM_data<=18'b100010110110011100;
        10'b1111011111:ROM_data<=18'b101101111011010001;
        10'b1111100000:ROM_data<=18'b011111111000000000;
        10'b1111100001:ROM_data<=18'b011110100110111000;
        10'b1111100010:ROM_data<=18'b011010101101110101;
        10'b1111100011:ROM_data<=18'b010100101100111110;
        10'b1111100100:ROM_data<=18'b011111111000000000;
        10'b1111100101:ROM_data<=18'b011000110101100000;
        10'b1111100110:ROM_data<=18'b000110100100000111;
        10'b1111100111:ROM_data<=18'b110001100100011101;
        10'b1111101000:ROM_data<=18'b011111111000000000;
        10'b1111101001:ROM_data<=18'b001111001100100000;
        10'b1111101010:ROM_data<=18'b101110101100101011;
        10'b1111101011:ROM_data<=18'b100000010000010100;
        10'b1111101100:ROM_data<=18'b011111111000000000;
        10'b1111101101:ROM_data<=18'b000011010100000011;
        10'b1111101110:ROM_data<=18'b100000111111001100;
        10'b1111101111:ROM_data<=18'b110110010011110010;
        10'b1111110000:ROM_data<=18'b011111111000000000;
        10'b1111110001:ROM_data<=18'b011101100110100000;
        10'b1111110010:ROM_data<=18'b010110110101001110;
        10'b1111110011:ROM_data<=18'b001100101100010111;
        10'b1111110100:ROM_data<=18'b011111111000000000;
        10'b1111110101:ROM_data<=18'b010110101101001101;
        10'b1111110110:ROM_data<=18'b000000011100000010;
        10'b1111110111:ROM_data<=18'b101010000101001001;
        10'b1111111000:ROM_data<=18'b011111111000000000;
        10'b1111111001:ROM_data<=18'b001100011100010110;
        10'b1111111010:ROM_data<=18'b101001110101001010;
        10'b1111111011:ROM_data<=18'b100010011001011101;
        10'b1111111100:ROM_data<=18'b011111111000000000;
        10'b1111111101:ROM_data<=18'b000000001100000010;
        10'b1111111110:ROM_data<=18'b100000010111111101;
        10'b1111111111:ROM_data<=18'b111111100011111110;

    endcase
  end
endmodule