
`resetall
`timescale 1ns/1ps
module ROM4_omega (ROM_data, ROM_addr,clk);
  
  parameter WORDLENGTH=18,ADDRLENGTH=8;
  
  output [WORDLENGTH-1:0] ROM_data;
  input 	[ADDRLENGTH-1:0] ROM_addr;
  input  clk;
  reg    [WORDLENGTH-1:0] ROM_data;


  always @ (posedge clk)
  begin
  case(ROM_addr)
8'b00000000:ROM_data<=18'b011111111000000000;
8'b00000001:ROM_data<=18'b011111111000000000;
8'b00000010:ROM_data<=18'b011111111000000000;
8'b00000011:ROM_data<=18'b011111111000000000;
8'b00000100:ROM_data<=18'b011111111000000000;
8'b00000101:ROM_data<=18'b011101011110011111;
8'b00000110:ROM_data<=18'b010110100101001100;
8'b00000111:ROM_data<=18'b001100001100010101;
8'b00001000:ROM_data<=18'b011111111000000000;
8'b00001001:ROM_data<=18'b010110100101001100;
8'b00001010:ROM_data<=18'b000000000100000001;
8'b00001011:ROM_data<=18'b101001100101001100;
8'b00001100:ROM_data<=18'b011111111000000000;
8'b00001101:ROM_data<=18'b001100001100010101;
8'b00001110:ROM_data<=18'b101001100101001100;
8'b00001111:ROM_data<=18'b100010101001100001;
8'b00010000:ROM_data<=18'b011111111000000000;
8'b00010001:ROM_data<=18'b011111101111101000;
8'b00010010:ROM_data<=18'b011111010111001111;
8'b00010011:ROM_data<=18'b011110100110110110;
8'b00010100:ROM_data<=18'b011111111000000000;
8'b00010101:ROM_data<=18'b011100000110001000;
8'b00010110:ROM_data<=18'b010001101100101100;
8'b00010111:ROM_data<=18'b000011000100000011;
8'b00011000:ROM_data<=18'b011111111000000000;
8'b00011001:ROM_data<=18'b010100001100111011;
8'b00011010:ROM_data<=18'b111001111100000110;
8'b00011011:ROM_data<=18'b100100000110001000;
8'b00011100:ROM_data<=18'b011111111000000000;
8'b00011101:ROM_data<=18'b001001010100001100;
8'b00011110:ROM_data<=18'b100101100101110011;
8'b00011111:ROM_data<=18'b100111011010100001;
8'b00100000:ROM_data<=18'b011111111000000000;
8'b00100001:ROM_data<=18'b011111010111001111;
8'b00100010:ROM_data<=18'b011101011110011111;
8'b00100011:ROM_data<=18'b011010100101110011;
8'b00100100:ROM_data<=18'b011111111000000000;
8'b00100101:ROM_data<=18'b011010100101110011;
8'b00100110:ROM_data<=18'b001100001100010101;
8'b00100111:ROM_data<=18'b111001111100000110;
8'b00101000:ROM_data<=18'b011111111000000000;
8'b00101001:ROM_data<=18'b010001101100101100;
8'b00101010:ROM_data<=18'b110011111100010101;
8'b00101011:ROM_data<=18'b100000110111001111;
8'b00101100:ROM_data<=18'b011111111000000000;
8'b00101101:ROM_data<=18'b000110001100000110;
8'b00101110:ROM_data<=18'b100010101110011111;
8'b00101111:ROM_data<=18'b101110011011010100;
8'b00110000:ROM_data<=18'b011111111000000000;
8'b00110001:ROM_data<=18'b011110100110110110;
8'b00110010:ROM_data<=18'b011010100101110011;
8'b00110011:ROM_data<=18'b010100001100111011;
8'b00110100:ROM_data<=18'b011111111000000000;
8'b00110101:ROM_data<=18'b011000101101011111;
8'b00110110:ROM_data<=18'b000110001100000110;
8'b00110111:ROM_data<=18'b110001000100100000;
8'b00111000:ROM_data<=18'b011111111000000000;
8'b00111001:ROM_data<=18'b001111000100100000;
8'b00111010:ROM_data<=18'b101110011100101100;
8'b00111011:ROM_data<=18'b100000011000011000;
8'b00111100:ROM_data<=18'b011111111000000000;
8'b00111101:ROM_data<=18'b000011000100000011;
8'b00111110:ROM_data<=18'b100000110111001111;
8'b00111111:ROM_data<=18'b110110110011110100;
8'b01000000:ROM_data<=18'b011111111000000000;
8'b01000001:ROM_data<=18'b011111110111111010;
8'b01000010:ROM_data<=18'b011111110111110100;
8'b01000011:ROM_data<=18'b011111110111101110;
8'b01000100:ROM_data<=18'b011111111000000000;
8'b01000101:ROM_data<=18'b011101001110011001;
8'b01000110:ROM_data<=18'b010101011101000100;
8'b01000111:ROM_data<=18'b001001111100001110;
8'b01001000:ROM_data<=18'b011111111000000000;
8'b01001001:ROM_data<=18'b010101111101001000;
8'b01001010:ROM_data<=18'b111110100100000010;
8'b01001011:ROM_data<=18'b100111111101011010;
8'b01001100:ROM_data<=18'b011111111000000000;
8'b01001101:ROM_data<=18'b001011011100010011;
8'b01001110:ROM_data<=18'b101000100101010101;
8'b01001111:ROM_data<=18'b100011101001110010;
8'b01010000:ROM_data<=18'b011111111000000000;
8'b01010001:ROM_data<=18'b011111101111100001;
8'b01010010:ROM_data<=18'b011110111111000011;
8'b01010011:ROM_data<=18'b011101101110100101;
8'b01010100:ROM_data<=18'b011111111000000000;
8'b01010101:ROM_data<=18'b011011101110000011;
8'b01010110:ROM_data<=18'b010000011100100110;
8'b01010111:ROM_data<=18'b000000110100000010;
8'b01011000:ROM_data<=18'b011111111000000000;
8'b01011001:ROM_data<=18'b010011100100110111;
8'b01011010:ROM_data<=18'b111000011100001001;
8'b01011011:ROM_data<=18'b100010111110011001;
8'b01011100:ROM_data<=18'b011111111000000000;
8'b01011101:ROM_data<=18'b001000100100001011;
8'b01011110:ROM_data<=18'b100100110101111101;
8'b01011111:ROM_data<=18'b101001000010101111;
8'b01100000:ROM_data<=18'b011111111000000000;
8'b01100001:ROM_data<=18'b011111000111001001;
8'b01100010:ROM_data<=18'b011100110110010011;
8'b01100011:ROM_data<=18'b011001001101100100;
8'b01100100:ROM_data<=18'b011111111000000000;
8'b01100101:ROM_data<=18'b011010000101101110;
8'b01100110:ROM_data<=18'b001010101100010000;
8'b01100111:ROM_data<=18'b110111100100001011;
8'b01101000:ROM_data<=18'b011111111000000000;
8'b01101001:ROM_data<=18'b010001000100101001;
8'b01101010:ROM_data<=18'b110010011100011010;
8'b01101011:ROM_data<=18'b100000011111100001;
8'b01101100:ROM_data<=18'b011111111000000000;
8'b01101101:ROM_data<=18'b000101011100000101;
8'b01101110:ROM_data<=18'b100010000110101011;
8'b01101111:ROM_data<=18'b110000011011011101;
8'b01110000:ROM_data<=18'b011111111000000000;
8'b01110001:ROM_data<=18'b011110010110110001;
8'b01110010:ROM_data<=18'b011001100101101001;
8'b01110011:ROM_data<=18'b010010010100110000;
8'b01110100:ROM_data<=18'b011111111000000000;
8'b01110101:ROM_data<=18'b011000001101011010;
8'b01110110:ROM_data<=18'b000100101100000100;
8'b01110111:ROM_data<=18'b101111000100101001;
8'b01111000:ROM_data<=18'b011111111000000000;
8'b01111001:ROM_data<=18'b001110010100011101;
8'b01111010:ROM_data<=18'b101101001100110100;
8'b01111011:ROM_data<=18'b100000101000101011;
8'b01111100:ROM_data<=18'b011111111000000000;
8'b01111101:ROM_data<=18'b000010010100000010;
8'b01111110:ROM_data<=18'b100000100111011011;
8'b01111111:ROM_data<=18'b111001001011111000;
8'b10000000:ROM_data<=18'b011111111000000000;
8'b10000001:ROM_data<=18'b011111110111110100;
8'b10000010:ROM_data<=18'b011111101111101000;
8'b10000011:ROM_data<=18'b011111100111011011;
8'b10000100:ROM_data<=18'b011111111000000000;
8'b10000101:ROM_data<=18'b011100110110010011;
8'b10000110:ROM_data<=18'b010100001100111011;
8'b10000111:ROM_data<=18'b000111101100001001;
8'b10001000:ROM_data<=18'b011111111000000000;
8'b10001001:ROM_data<=18'b010101011101000100;
8'b10001010:ROM_data<=18'b111101000100000011;
8'b10001011:ROM_data<=18'b100110100101101001;
8'b10001100:ROM_data<=18'b011111111000000000;
8'b10001101:ROM_data<=18'b001010101100010000;
8'b10001110:ROM_data<=18'b100111011101011111;
8'b10001111:ROM_data<=18'b100100110010000011;
8'b10010000:ROM_data<=18'b011111111000000000;
8'b10010001:ROM_data<=18'b011111100111011011;
8'b10010010:ROM_data<=18'b011110100110110110;
8'b10010011:ROM_data<=18'b011100110110010011;
8'b10010100:ROM_data<=18'b011111111000000000;
8'b10010101:ROM_data<=18'b011011010101111101;
8'b10010110:ROM_data<=18'b001111000100100000;
8'b10010111:ROM_data<=18'b111110100100000010;
8'b10011000:ROM_data<=18'b011111111000000000;
8'b10011001:ROM_data<=18'b010010111100110100;
8'b10011010:ROM_data<=18'b110110110100001100;
8'b10011011:ROM_data<=18'b100010000110101011;
8'b10011100:ROM_data<=18'b011111111000000000;
8'b10011101:ROM_data<=18'b000111101100001001;
8'b10011110:ROM_data<=18'b100100000110001000;
8'b10011111:ROM_data<=18'b101010101010111100;
8'b10100000:ROM_data<=18'b011111111000000000;
8'b10100001:ROM_data<=18'b011110111111000011;
8'b10100010:ROM_data<=18'b011100000110001000;
8'b10100011:ROM_data<=18'b010111100101010101;
8'b10100100:ROM_data<=18'b011111111000000000;
8'b10100101:ROM_data<=18'b011001100101101001;
8'b10100110:ROM_data<=18'b001001010100001100;
8'b10100111:ROM_data<=18'b110101011100010000;
8'b10101000:ROM_data<=18'b011111111000000000;
8'b10101001:ROM_data<=18'b010000011100100110;
8'b10101010:ROM_data<=18'b110001000100100000;
8'b10101011:ROM_data<=18'b100000010111110100;
8'b10101100:ROM_data<=18'b011111111000000000;
8'b10101101:ROM_data<=18'b000100101100000100;
8'b10101110:ROM_data<=18'b100001100110110110;
8'b10101111:ROM_data<=18'b110010011011100110;
8'b10110000:ROM_data<=18'b011111111000000000;
8'b10110001:ROM_data<=18'b011110000110101011;
8'b10110010:ROM_data<=18'b011000101101011111;
8'b10110011:ROM_data<=18'b010000011100100110;
8'b10110100:ROM_data<=18'b011111111000000000;
8'b10110101:ROM_data<=18'b010111100101010101;
8'b10110110:ROM_data<=18'b000011000100000011;
8'b10110111:ROM_data<=18'b101101001100110100;
8'b10111000:ROM_data<=18'b011111111000000000;
8'b10111001:ROM_data<=18'b001101101100011010;
8'b10111010:ROM_data<=18'b101011111100111011;
8'b10111011:ROM_data<=18'b100001001000111101;
8'b10111100:ROM_data<=18'b011111111000000000;
8'b10111101:ROM_data<=18'b000001100100000010;
8'b10111110:ROM_data<=18'b100000011111101000;
8'b10111111:ROM_data<=18'b111011011011111100;
8'b11000000:ROM_data<=18'b011111111000000000;
8'b11000001:ROM_data<=18'b011111110111101110;
8'b11000010:ROM_data<=18'b011111100111011011;
8'b11000011:ROM_data<=18'b011111000111001001;
8'b11000100:ROM_data<=18'b011111111000000000;
8'b11000101:ROM_data<=18'b011100011110001110;
8'b11000110:ROM_data<=18'b010010111100110100;
8'b11000111:ROM_data<=18'b000101011100000101;
8'b11001000:ROM_data<=18'b011111111000000000;
8'b11001001:ROM_data<=18'b010100110100111111;
8'b11001010:ROM_data<=18'b111011011100000100;
8'b11001011:ROM_data<=18'b100101001101111000;
8'b11001100:ROM_data<=18'b011111111000000000;
8'b11001101:ROM_data<=18'b001001111100001110;
8'b11001110:ROM_data<=18'b100110100101101001;
8'b11001111:ROM_data<=18'b100110000010010010;
8'b11010000:ROM_data<=18'b011111111000000000;
8'b11010001:ROM_data<=18'b011111011111010101;
8'b11010010:ROM_data<=18'b011110000110101011;
8'b11010011:ROM_data<=18'b011011101110000011;
8'b11010100:ROM_data<=18'b011111111000000000;
8'b11010101:ROM_data<=18'b011010111101111000;
8'b11010110:ROM_data<=18'b001101101100011010;
8'b11010111:ROM_data<=18'b111100001100000011;
8'b11011000:ROM_data<=18'b011111111000000000;
8'b11011001:ROM_data<=18'b010010010100110000;
8'b11011010:ROM_data<=18'b110101011100010000;
8'b11011011:ROM_data<=18'b100001011110111100;
8'b11011100:ROM_data<=18'b011111111000000000;
8'b11011101:ROM_data<=18'b000110111100001000;
8'b11011110:ROM_data<=18'b100011010110010011;
8'b11011111:ROM_data<=18'b101100100011001001;
8'b11100000:ROM_data<=18'b011111111000000000;
8'b11100001:ROM_data<=18'b011110101110111100;
8'b11100010:ROM_data<=18'b011011010101111101;
8'b11100011:ROM_data<=18'b010101111101001000;
8'b11100100:ROM_data<=18'b011111111000000000;
8'b11100101:ROM_data<=18'b011001001101100100;
8'b11100110:ROM_data<=18'b000111101100001001;
8'b11100111:ROM_data<=18'b110011001100010111;
8'b11101000:ROM_data<=18'b011111111000000000;
8'b11101001:ROM_data<=18'b001111101100100011;
8'b11101010:ROM_data<=18'b101111101100100110;
8'b11101011:ROM_data<=18'b100000010000000110;
8'b11101100:ROM_data<=18'b011111111000000000;
8'b11101101:ROM_data<=18'b000011111100000011;
8'b11101110:ROM_data<=18'b100001001111000011;
8'b11101111:ROM_data<=18'b110100101011101101;
8'b11110000:ROM_data<=18'b011111111000000000;
8'b11110001:ROM_data<=18'b011101101110100101;
8'b11110010:ROM_data<=18'b010111100101010101;
8'b11110011:ROM_data<=18'b001110010100011101;
8'b11110100:ROM_data<=18'b011111111000000000;
8'b11110101:ROM_data<=18'b010111000101010001;
8'b11110110:ROM_data<=18'b000001100100000010;
8'b11110111:ROM_data<=18'b101011010100111111;
8'b11111000:ROM_data<=18'b011111111000000000;
8'b11111001:ROM_data<=18'b001100111100010111;
8'b11111010:ROM_data<=18'b101010101101000100;
8'b11111011:ROM_data<=18'b100001110001001111;
8'b11111100:ROM_data<=18'b011111111000000000;
8'b11111101:ROM_data<=18'b000000110100000010;
8'b11111110:ROM_data<=18'b100000010111110100;
8'b11111111:ROM_data<=18'b111101110011111110;
  endcase

//    ROM_data<=ROM[ROM_addr];
  end
  
  
//  initial $readmemb ("w_im_bin_flow4.txt",  ROM);
endmodule