
//
// using Mentor Graphics HDL Designer(TM) 2004.1b (Build 12)
//
`resetall
`timescale 1ns/1ps
module ROM3_omega (ROM_data, ROM_addr,clk);
  
  parameter WORDLENGTH=18,ADDRLENGTH=6;
  
  output [WORDLENGTH-1:0] ROM_data;
  input 	[ADDRLENGTH-1:0] ROM_addr;
  input  clk;
  reg    [WORDLENGTH-1:0] ROM_data;
  
  always @ (posedge clk)
  begin
    case(ROM_addr)
6'b000000:ROM_data<=18'b011111111000000000;
6'b000001:ROM_data<=18'b011111111000000000;
6'b000010:ROM_data<=18'b011111111000000000;
6'b000011:ROM_data<=18'b011111111000000000;
6'b000100:ROM_data<=18'b011111111000000000;
6'b000101:ROM_data<=18'b011101011110011111;
6'b000110:ROM_data<=18'b010110100101001100;
6'b000111:ROM_data<=18'b001100001100010101;
6'b001000:ROM_data<=18'b011111111000000000;
6'b001001:ROM_data<=18'b010110100101001100;
6'b001010:ROM_data<=18'b000000000100000001;
6'b001011:ROM_data<=18'b101001100101001100;
6'b001100:ROM_data<=18'b011111111000000000;
6'b001101:ROM_data<=18'b001100001100010101;
6'b001110:ROM_data<=18'b101001100101001100;
6'b001111:ROM_data<=18'b100010101001100001;
6'b010000:ROM_data<=18'b011111111000000000;
6'b010001:ROM_data<=18'b011111101111101000;
6'b010010:ROM_data<=18'b011111010111001111;
6'b010011:ROM_data<=18'b011110100110110110;
6'b010100:ROM_data<=18'b011111111000000000;
6'b010101:ROM_data<=18'b011100000110001000;
6'b010110:ROM_data<=18'b010001101100101100;
6'b010111:ROM_data<=18'b000011000100000011;
6'b011000:ROM_data<=18'b011111111000000000;
6'b011001:ROM_data<=18'b010100001100111011;
6'b011010:ROM_data<=18'b111001111100000110;
6'b011011:ROM_data<=18'b100100000110001000;
6'b011100:ROM_data<=18'b011111111000000000;
6'b011101:ROM_data<=18'b001001010100001100;
6'b011110:ROM_data<=18'b100101100101110011;
6'b011111:ROM_data<=18'b100111011010100001;
6'b100000:ROM_data<=18'b011111111000000000;
6'b100001:ROM_data<=18'b011111010111001111;
6'b100010:ROM_data<=18'b011101011110011111;
6'b100011:ROM_data<=18'b011010100101110011;
6'b100100:ROM_data<=18'b011111111000000000;
6'b100101:ROM_data<=18'b011010100101110011;
6'b100110:ROM_data<=18'b001100001100010101;
6'b100111:ROM_data<=18'b111001111100000110;
6'b101000:ROM_data<=18'b011111111000000000;
6'b101001:ROM_data<=18'b010001101100101100;
6'b101010:ROM_data<=18'b110011111100010101;
6'b101011:ROM_data<=18'b100000110111001111;
6'b101100:ROM_data<=18'b011111111000000000;
6'b101101:ROM_data<=18'b000110001100000110;
6'b101110:ROM_data<=18'b100010101110011111;
6'b101111:ROM_data<=18'b101110011011010100;
6'b110000:ROM_data<=18'b011111111000000000;
6'b110001:ROM_data<=18'b011110100110110110;
6'b110010:ROM_data<=18'b011010100101110011;
6'b110011:ROM_data<=18'b010100001100111011;
6'b110100:ROM_data<=18'b011111111000000000;
6'b110101:ROM_data<=18'b011000101101011111;
6'b110110:ROM_data<=18'b000110001100000110;
6'b110111:ROM_data<=18'b110001000100100000;
6'b111000:ROM_data<=18'b011111111000000000;
6'b111001:ROM_data<=18'b001111000100100000;
6'b111010:ROM_data<=18'b101110011100101100;
6'b111011:ROM_data<=18'b100000011000011000;
6'b111100:ROM_data<=18'b011111111000000000;
6'b111101:ROM_data<=18'b000011000100000011;
6'b111110:ROM_data<=18'b100000110111001111;
6'b111111:ROM_data<=18'b110110110011110100;

    endcase
  end
endmodule